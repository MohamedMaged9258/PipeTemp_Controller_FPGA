library verilog;
use verilog.vl_types.all;
entity PipeTemp_Controller_tb is
end PipeTemp_Controller_tb;
